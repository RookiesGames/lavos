module plugins

enum Platform {
	android
	ios
}
